** Generated for: hspiceD
** Generated on: Nov  9 17:26:08 2022
** Design library name: cad3
** Design cell name: loaded_nand
** Design view name: schematic
.GLOBAL vss! vdd!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad3
** Cell name: NAND2
** View name: schematic
*.subckt NAND2 a b z
*mnmos1 net1 b vss! vss! NMOS_VTL L=50e-9 W=300e-9 AD=31.5e-15 AS=31.5e-15 PD=510e-9 PS=510e-9 M=1
*mnmos0 z a net1 vss! NMOS_VTL L=50e-9 W=300e-9 AD=31.5e-15 AS=31.5e-15 PD=510e-9 PS=510e-9 M=1
*mpmos0 z a vdd! vdd! PMOS_VTL L=50e-9 W=250e-9 AD=26.25e-15 AS=26.25e-15 PD=460e-9 PS=460e-9 M=1
*mpmos1 z b vdd! vdd! PMOS_VTL L=50e-9 W=250e-9 AD=26.25e-15 AS=26.25e-15 PD=460e-9 PS=460e-9 M=1
*.ends NAND2
** End of subcircuit definition.

** ==== Post - layout netlist ====
.include loaded_nand.pex.netlist

** ==== loaded_inverter circuit ====
** Library name: cad3
** Cell name: loaded_nand
** View name: schematic
xdut a b z NAND2
xnand3 vdd! z net5 NAND2
xnand2 vdd! z net4 NAND2
xnand1 vdd! z net2 NAND2
xnand0 vdd! z net3 NAND2
.END
