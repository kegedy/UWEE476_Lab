.GLOBAL vdd!


.OPTION

m0 vo vi 0 0 NMOS_VTL L=50e-9 W=1e-6 AD=105e-15 AS=105e-15 PD=1.21e-6 PS=1.21e-6 M=1
r0 vdd! vo 100e3
.END
