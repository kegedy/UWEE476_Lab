** Generated for: hspiceD
** Generated on: Oct 21 19:00:39 2022
** Design library name: cad1
** Design cell name: q4
** Design view name: schematic
.GLOBAL vdd!


.TEMP 25
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad1
** Cell name: q4
** View name: schematic
m0 vdd! vin vdd! vdd! NMOS_VTL L=50e-9 W=1e-6 AD=105e-15 AS=105e-15 PD=1.21e-6 PS=1.21e-6 M=1
.END
