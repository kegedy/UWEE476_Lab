* SPICE NETLIST
***************************************

.SUBCKT AlphaPhaseLatch Clk_rst Q Q_bar rst D Clk VSS! VDD!
** N=17 EP=8 IP=0 FDC=22
M0 Q Clk_rst Q VSS! NMOS_VTL L=1.65e-07 W=1.5e-07 AD=2.325e-14 AS=2.325e-14 PD=4.55e-07 PS=4.55e-07 $X=255 $Y=905 $D=1
M1 3 Clk Q VSS! NMOS_VTL L=5e-08 W=3e-07 AD=3.15e-14 AS=4.65e-14 PD=8.1e-07 PS=9.1e-07 $X=425 $Y=905 $D=1
M2 VSS! Q Q_bar VSS! NMOS_VTL L=5e-08 W=3e-07 AD=4.35e-14 AS=4.65e-14 PD=8.9e-07 PS=9.1e-07 $X=815 $Y=905 $D=1
M3 6 Q_bar VSS! VSS! NMOS_VTL L=5e-08 W=3e-07 AD=4.35e-14 AS=4.35e-14 PD=8.9e-07 PS=8.9e-07 $X=1010 $Y=905 $D=1
M4 VSS! rst 6 VSS! NMOS_VTL L=5e-08 W=3e-07 AD=3.15e-14 AS=4.35e-14 PD=8.1e-07 PS=8.9e-07 $X=1205 $Y=905 $D=1
M5 7 Q_bar VSS! VSS! NMOS_VTL L=5e-08 W=3e-07 AD=4.35e-14 AS=3.15e-14 PD=8.9e-07 PS=8.1e-07 $X=1545 $Y=905 $D=1
M6 VSS! 6 7 VSS! NMOS_VTL L=5e-08 W=3e-07 AD=4.35e-14 AS=4.35e-14 PD=8.9e-07 PS=8.9e-07 $X=1740 $Y=905 $D=1
M7 8 6 VSS! VSS! NMOS_VTL L=5e-08 W=3e-07 AD=4.35e-14 AS=4.35e-14 PD=8.9e-07 PS=8.9e-07 $X=1935 $Y=905 $D=1
M8 VSS! rst 8 VSS! NMOS_VTL L=5e-08 W=3e-07 AD=3.15e-14 AS=4.35e-14 PD=8.1e-07 PS=8.9e-07 $X=2130 $Y=905 $D=1
M9 3 8 VSS! VSS! NMOS_VTL L=5e-08 W=3e-07 AD=4.35e-14 AS=3.15e-14 PD=8.9e-07 PS=8.1e-07 $X=2470 $Y=905 $D=1
M10 VSS! 7 3 VSS! NMOS_VTL L=5e-08 W=3e-07 AD=3.15e-14 AS=4.35e-14 PD=8.1e-07 PS=8.9e-07 $X=2665 $Y=905 $D=1
M11 Q Clk D VDD! PMOS_VTL L=5e-08 W=4e-07 AD=6.2e-14 AS=4.2e-14 PD=1.11e-06 PS=1.01e-06 $X=220 $Y=1515 $D=0
M12 3 Clk_rst Q VDD! PMOS_VTL L=5e-08 W=4e-07 AD=4.2e-14 AS=6.2e-14 PD=1.01e-06 PS=1.11e-06 $X=425 $Y=1515 $D=0
M13 VDD! Q Q_bar VDD! PMOS_VTL L=5e-08 W=4e-07 AD=5.8e-14 AS=6.2e-14 PD=1.09e-06 PS=1.11e-06 $X=815 $Y=1515 $D=0
M14 14 Q_bar VDD! VDD! PMOS_VTL L=5e-08 W=4e-07 AD=5.8e-14 AS=5.8e-14 PD=1.09e-06 PS=1.09e-06 $X=1010 $Y=1515 $D=0
M15 6 rst 14 VDD! PMOS_VTL L=5e-08 W=4e-07 AD=4.2e-14 AS=5.8e-14 PD=1.01e-06 PS=1.09e-06 $X=1205 $Y=1515 $D=0
M16 15 Q_bar 7 VDD! PMOS_VTL L=5e-08 W=4e-07 AD=5.8e-14 AS=4.2e-14 PD=1.09e-06 PS=1.01e-06 $X=1545 $Y=1515 $D=0
M17 VDD! 6 15 VDD! PMOS_VTL L=5e-08 W=4e-07 AD=5.8e-14 AS=5.8e-14 PD=1.09e-06 PS=1.09e-06 $X=1740 $Y=1515 $D=0
M18 16 6 VDD! VDD! PMOS_VTL L=5e-08 W=4e-07 AD=5.8e-14 AS=5.8e-14 PD=1.09e-06 PS=1.09e-06 $X=1935 $Y=1515 $D=0
M19 8 rst 16 VDD! PMOS_VTL L=5e-08 W=4e-07 AD=4.2e-14 AS=5.8e-14 PD=1.01e-06 PS=1.09e-06 $X=2130 $Y=1515 $D=0
M20 17 8 3 VDD! PMOS_VTL L=5e-08 W=4e-07 AD=5.8e-14 AS=4.2e-14 PD=1.09e-06 PS=1.01e-06 $X=2470 $Y=1515 $D=0
M21 VDD! 7 17 VDD! PMOS_VTL L=5e-08 W=4e-07 AD=4.2e-14 AS=5.8e-14 PD=1.01e-06 PS=1.09e-06 $X=2665 $Y=1515 $D=0
.ENDS
***************************************
