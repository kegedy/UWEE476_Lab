** Generated for: hspiceD
** Generated on: Oct 14 17:20:10 2022
** Design library name: cad1
** Design cell name: q1d_1
** Design view name: schematic
.GLOBAL vdd!
.PARAM vdrain


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad1
** Cell name: q1d_1
** View name: schematic
m0 net1 vin vdd! vdd! PMOS_VTL L=50e-9 W=1e-6 AD=105e-15 AS=105e-15 PD=1.21e-6 PS=1.21e-6 M=1
v0 net1 0 DC=vdrain
.END
