** Generated for: hspiceD
** Generated on: Nov 14 05:39:02 2022
** Design library name: cad3
** Design cell name: NAND2_balanced
** Design view name: schematic
.GLOBAL vdd! vss!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad3
** Cell name: NAND2_balanced
** View name: schematic
mnmos1 net1 b vss! vss! NMOS_VTL L=50e-9 W=300e-9 AD=31.5e-15 AS=31.5e-15 PD=510e-9 PS=510e-9 M=1
mnmos0 out a net1 vss! NMOS_VTL L=50e-9 W=300e-9 AD=31.5e-15 AS=31.5e-15 PD=510e-9 PS=510e-9 M=1
mpmos0 out a vdd! vdd! PMOS_VTL L=50e-9 W=250e-9 AD=26.25e-15 AS=26.25e-15 PD=460e-9 PS=460e-9 M=1
mpmos1 out b vdd! vdd! PMOS_VTL L=50e-9 W=250e-9 AD=26.25e-15 AS=26.25e-15 PD=460e-9 PS=460e-9 M=1
.END
