** Generated for: hspiceD
** Generated on: Oct 14 14:31:22 2022
** Design library name: cad1
** Design cell name: q1c
** Design view name: schematic
.GLOBAL vdd!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad1
** Cell name: q1c
** View name: schematic
m0 0 vin vdd! vdd! PMOS_VTL L=50e-9 W=1e-6 AD=105e-15 AS=105e-15 PD=1.21e-6 PS=1.21e-6 M=1
.END
