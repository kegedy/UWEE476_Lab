../netlists/nmos_inverter/hspiceD/schematic/netlist/input.ckt