** Generated for: hspiceD
** Generated on: Oct 14 13:19:33 2022
** Design library name: cad1
** Design cell name: q1b_2
** Design view name: schematic
.GLOBAL vdd!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad1
** Cell name: q1b_2
** View name: schematic
m0 vdd! vin 0 0 NMOS_VTL L=50e-9 W=1e-6 AD=105e-15 AS=105e-15 PD=1.21e-6 PS=1.21e-6 M=1
.END
