../netlists/rc_series/hspiceD/schematic/netlist/input.ckt