** Generated for: hspiceD
** Generated on: Oct 14 19:34:58 2022
** Design library name: cad1
** Design cell name: q2a_2
** Design view name: schematic
.GLOBAL vdd!


.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2

** Library name: cad1
** Cell name: q2a_2
** View name: schematic
m0 vo vi 0 0 NMOS_VTL L=50e-9 W=1e-6 AD=105e-15 AS=105e-15 PD=1.21e-6 PS=1.21e-6 M=1
r0 vdd! vo 200e3
.END
